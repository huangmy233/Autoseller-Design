`timescale 1ns/1ps
module Autoseller_tb2;